module note_gen(
    clk, // clock from crystal
    rst, // active high reset
    // volume, 
    // note_div_left, // div for note generation
    note_div,
    // audio_left,
    audio
);

    // I/O declaration
    input clk; // clock from crystal
    input rst; // active low reset
    // input [2:0] volume;
    input [21:0] note_div; // div for note generation
    output [15:0] audio;

    // Declare internal signals
    reg [21:0] clk_cnt_next, clk_cnt;
    reg [21:0] clk_cnt_next_2, clk_cnt_2;
    reg b_clk, b_clk_next;
    reg c_clk, c_clk_next;

    // Note frequency generation
    // clk_cnt, clk_cnt_2, b_clk, c_clk
    always @(posedge clk or posedge rst)
        if (rst == 1'b1)
            begin
                // clk_cnt <= 22'd0;
                clk_cnt_2 <= 22'd0;
                // b_clk <= 1'b0;
                c_clk <= 1'b0;
            end
        else
            begin
                // clk_cnt <= clk_cnt_next;
                clk_cnt_2 <= clk_cnt_next_2;
                // b_clk <= b_clk_next;
                c_clk <= c_clk_next;
            end
    
    // clk_cnt_next, b_clk_next
    // always @*
    //     if (clk_cnt == note_div_left)
    //         begin
    //             clk_cnt_next = 22'd0;
    //             b_clk_next = ~b_clk;
    //         end
    //     else
    //         begin
    //             clk_cnt_next = clk_cnt + 1'b1;
    //             b_clk_next = b_clk;
    //         end

    // clk_cnt_next_2, c_clk_next
    always @*
        if (clk_cnt_2 == note_div)
            begin
                clk_cnt_next_2 = 22'd0;
                c_clk_next = ~c_clk;
            end
        else
            begin
                clk_cnt_next_2 = clk_cnt_2 + 1'b1;
                c_clk_next = c_clk;
            end

    // Assign the amplitude of the note
    // Volume is controlled here
    // assign audio_left = (note_div_left == 22'd1) ? 16'h0000 : 
    //                             (b_clk == 1'b0) ? 16'hE000 : 16'h2000;
    assign audio = (note_div == 22'd1) ? 16'h0000 : 
                                (c_clk == 1'b0) ? 16'hE000 : 16'h2000;
endmodule